b0VIM 7.2      ���Uҁ�
8E  w                                       localhost.localdomain                   ~w/huarzail/CMP_POPNET/program/allShortPath/cluster0/hello.c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 utf-8U3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           �                            j       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ad     �     �       �  �  �  �  �  �  �  �  k  P  5    �  �  �  �  �  �  w  \  A  &    �  �  �  �  �  �  �  �  n  O  -  ,  �  �  �  �  �  �  �  �  h  F  %        �  �  �  �  �  �  }  w  _  H  7    �
  �
  �
  �
  �
  f
  X
  7
  
  �	  �	  �	  �	  �	  }	  m	  R	  0	  	  	  �  �  �  �  �  v  k  <  &    �  �  �  �  }  {  z  U  J  1      �  �  �  �  �  �  ^  ;  5  4  2  1  $  �  �  �  �  �  X  Q  5    �  �  �  �  �  �  �  |  e  _  I  G  F        �  �  �  �  �  �  r  k  h  [  4         �  �  �  �  �  �  �  �          }     }         a[i]=b[i];     for(i=0;i<NODENUM;i++){     int i; void CopyArray(int a[NODENUM],int b[NODENUM]){  }     fflush(stdout);     printf("Write file is over...\n"); 	fclose(fp); 	} 		i++;         fprintf(fp,"%d ",array[i]); 	{ 	while(i<n) 	fp=fopen(contents,"w");     fflush(stdout);     printf("Write file is beginning...\n"); 	int i=0; 	FILE *fp; { void WriteFile(char *contents,int array[],int n)  }     dist[destNo] = 0;     }         dist[i] = INF;     for(i=0; i<NODENUM; i++){     int i; void InitialDist(int dist[NODENUM],int destNo){   }     MTA_printresult();     fflush(stdout);     printf("leaving MTA_acquiesce..........\n");     *receiveSignal0 = 0x55;     }	          MTA_acquiesce(receiveSignal0); 	while(0xaa != *receiveSignal0){     MTA_printresult();     fflush(stdout);     printf("entering MTA_acquiesce.......... \n"); 	int *receiveSignal0= (int *)cmp0_5; void Wait(){  }      } 	    dist[i] = *receiveAddress0++; 	for(i=LOCALNUM; i<NODENUM; i++){     int *receiveAddress0= (int *)cmp0_0; 	int i; void ReceiveData(int dist[NODENUM]){ }     fflush(stdout);         printf("\n");	         }             printf("%d\t",dist[i]); 	for(i=0;i<NODENUM;i++){     int i; void PrintResult(int dist[NODENUM]){  }     *(localAddress0+node) = tmp[node];     }         } 		    tmp[node]= c[node][i] + dist[i];          if(c[node][i]+dist[i] < tmp[node]){     for(i=0; i<NODENUM; i++){         tmp[i] = INF;     for(i=0;i<LOCALNUM;i++)//initial the tmp[]     int i;     int tmp[LOCALNUM]; 	int *localAddress0 = (int *)cmp0_2; void CulculateMin(int node, int dist[NODENUM], int c[NODENUM][NODENUM]){  }     }         }             if(i==j) c[i][j] = 0;         for(j=0; j<NODENUM; j++){ 	for(i=0; i<NODENUM; i++){     fclose(fp);     printf("\n");     }         c[a[1]][a[0]]=a[2];         c[a[0]][a[1]]=a[2];                 if(i == 3) i=0;                     printf("\n");                     printf("%d ",a[i]);                 for(i=0;i<3;i++)             }                 p=strtok(NULL," ");                 i++;                 a[i] = atoi(p);             {             while (p)             p=strtok(str," ");         if (fgets(str,sizeof(str),fp)==NULL) break ;         char *p;         memset(a,0,3);         char str[1024];     {     while(!feof(fp))         }         printf("open file error\n");     {     if (fp == NULL)     fp=fopen(contents,"r");     //begin to read file          }         }             else  c[i][j] = INF;             if(i==j) c[i][j] = 0;         for(j=0; j<NODENUM; j++){     for(i=0; i<NODENUM; i++){     //initialization      FILE *fp;     int a[3];     int j;     int i = 0; void ReadFile(char *contents, int c[NODENUM][NODENUM]){  volatile int x[NODENUM][NODENUM]; volatile int DistTmp[NODENUM]; volatile int Dist[NODENUM];  #define MULTIPLE 2 #define INITIALNUM 255 #define LOCALNUM 128 #define NODENUM 256 #define INF 9999  #define cmp1_7 0x1ff008000 #define cmp1_6 0x1ff007000 #define cmp1_5 0x1ff006000 #define cmp1_4 0x1ff005000 #define cmp1_3 0x1ff004000 #define cmp1_2 0x1ff003000 #define cmp1_1 0x1ff002000 #define cmp1_0 0x1ff001000  #define cmp0_6 0x11fde6f50 #define cmp0_5 0x1ff000800 #define cmp0_4 0x1ff000400 #define cmp0_3 0x1ff000300 #define cmp0_2 0x1ff000200 #define cmp0_1 0x1ff000100 #define cmp0_0 0x1ff000000  volatile int CountLock = 0; #define NPROC 64  #include "stdint.h" #include "barrier.h" #include "stdio.h" #define global ad  e  )     j       �  �  �  �  �  �  �  e  I  %  �  �  �  �  �  �  �  l  P  J  *  #    �  �  �  �  l  ,      �  �  �  �  �  �  �  �  a  G  F  3  
  �  �  �  �  _  ^  G  *  �
  �
  �
  �
  K
  
  �	  �	  �	  �	  �	  �	  �	  �	  Q	  P	  	  �    G  5  4     �  �  �  �  j  T  S  I  1  �  �  �  F  E  ;  #  �  �  �  �  �  �  ^  K  <  1  /  .  ,  +  )  -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	  	  } 	while(1); 	MTA_Stats(0); 	MTA_Bar_Stats(0); 	barrier(MTA_getthreadID() , NPROC); 	MTA_Bar_Stats(1); 	}         } 		    WriteFile("./output.txt",Dist,NODENUM);             PrintResult(Dist);             printf("The simulation result is:\n");         if(my_id == 0){         }              printf("****************print the final cycle end********************\n");             MTA_printresult();             fflush(stdout);             printf("****************print the final cycle begin********************\n");         if(my_id == 0){         }  			MTA_Bar_Stats(0);	 			barrier(MTA_getthreadID() , NPROC); 			MTA_Bar_Stats(1); 			}			                 fflush(stdout);                 printf("I received the data.\n"); 				ReceiveData(Dist);//receive the other Dist[]			  				Wait();//wait                 printf("Cluster0 sending is over!\n");  				//MTA_mailboxsend(0,localSignal0,1,otherSignal0,1,1);//send signal 				MTA_mailboxsend(0,localAddress2,1,otherAddress0,LOCALNUM,1);//send the data     				printf("Data from cluster0 send to cluster1.\n");                  CopyArray(Dist,DistTmp);                      if(my_id == 0){	  			MTA_Bar_Stats(0); 			barrier(MTA_getthreadID() , NPROC); 			MTA_Bar_Stats(1); 	                 } 		    DistTmp[MULTIPLE*my_id+i] = *(localAddress1+MULTIPLE*my_id+i); 			CulculateMin(MULTIPLE*my_id+i, Dist, x);//culculate the minimize			         for(i=0;i<MULTIPLE;i++){             }                 fflush(stdout);                 printf("**********This is the %dth loop**********\n",k);             if (my_id == 3){ 		for(k=0; k<80; k++){          int *localSignal0   =   (int *)cmp0_1;  		int *localAddress2  =   (int *)cmp0_2; 		int *localAddress1  =   (int *)cmp0_2; 		int *otherSignal0   =   (int *)cmp1_1; 		int *otherAddress0  =   (int *)cmp1_0;         int i,j,k;          //fflush(stdout); 		//printf("come on after fork %d.\n",my_id); 		my_id = MTA_getthreadID();  	{ 	MTA_Stats(1);  	MTA_Bar_Stats(0);	 	barrier(MTA_getthreadID() , NPROC); 	MTA_Bar_Stats(1); 	}     		if(my_id != 0)		break; 		printf("loop %d after MTA_getthreadID %d\n",ProcessId,my_id); 		my_id = MTA_getthreadID(); 		printf("loop %d after fork %d\n",ProcessId,my_id); 		my_id = MTA_fork();     { 	for(ProcessId = 1;ProcessId < NPROC; ProcessId++) 	barrier_init(NPROC);     }          printf("%d\t",Dist[i]);     {     for(i=0; i<NODENUM;i++)     printf("The orignal dist[] is:\n");         InitialDist(Dist,INITIALNUM);//initialization       }             printf("\n");             }                    printf("%d ", x[i][j]);             for(j=0;j<NODENUM;j++){     for(i=0;i<NODENUM;i++){     printf("The orignal x[][] is:\n");     ReadFile("./input.txt",x);//read file      int i,j,cnt=0; 	int my_id = 0; 	unsigned ProcessId = 0; { int main() 