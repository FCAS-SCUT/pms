b0VIM 7.3      ��]Uo�W!K  w                                       localhost.localdomain                   ~w/huarzail/CMP_POPNET/program/fastSort/cluster0/hello.c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     utf-8U3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           �                     ��������w       �                     0       "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     ad     �     �       �  �  �  �  �  �  �  �  k  P  5    �  �  �  �  �  �  w  \  A  &    �  �  �  �  �  �  �  �  �  p  J  I         �  �  �  �  �  �  |  v  ]  W  ?  .  �  �  �  �  �  �  ]  O  >  8  &        �
  �
  �
  �
  �
  |
  r
  g
  Y
  U
  4
  
  
  
  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  n	  k	  Y	  @	  	  	  	  �  �  �  �  �  �  �  �  z  n  j  g  T  G  &      �  �  �  �  j  V  7    �  �  �  t  K  2  0  /  
  �  �  �  �  �  �  �  h  `  7    �  �  �  �  �  �  �  �  x  d  K  ?         	  �  �  �  �  �  �  g  K  #        �  �  �             	int i; void InitialDist(int coreNum,int array[],int x[],int *p, int *q){  }     }	          MTA_acquiesce(receiveSignal0); 	while(*receiveSignal0!=a){     *receiveSignal0 = 0;//receive signal 	int *receiveSignal0= (int *)cmp0_5; void WaitTime(int a){  }     fflush(stdout);     printf("Write file is over...\n"); 	fclose(fp); 	} 		i++; 		{fprintf(fp,"%d ",array[i]); 	while(i<n) 	fp=fopen(contents,"w");     fflush(stdout);     printf("Write file is beginning...\n"); 	int i=0; 	FILE *fp; { void WriteFile(char *contents,int array[],int n)  }     } 	    c[i] = *receiveAddress0++; 	for(i=LOCALNUM; i<NODENUM; i++){     int *receiveAddress0= (int *)cmp0_0; 	int i; void ReceiveData(int c[NODENUM]){ }     fflush(stdout);         printf("\n");	         }             printf("%d ",dist[i]); 	for(i=0;i<NODENUM+2;i++){     int i; void PrintResult(int dist[NODENUM]){  } 		arr[i] = newarr[p];    	for(i=low,p=0;p<(high-low+1);i++,p++)   	while(j<=high)     newarr[p++] = arr[j++];      	while(i<=mid)     newarr[p++] = arr[i++];    	}      		else      newarr[p++] = arr[j++];    		if(arr[i] < arr[j])   newarr[p++] = arr[i++];      	while(i<=mid && j<=high){         fflush(stdout);     printf("The merge_sort is beginning...\n"); 	int newarr[100000]; 	int i=low,j=mid+1,p=0;    {  void MergeSort(int arr[],int low,int mid, int high) }      QuickSortSecond(i+1,right,a);     QuickSortSecond(left,i-1,a); 	a[i]=temp;      a[left]=a[i];  	} 		} 			a[j]=t;  			a[i]=a[j];  			t=a[i];  		{  		if(i<j)  		while(a[i]<=temp && i<j) i++;  		while(a[j]>=temp && i<j) j--;  	{  	while(i!=j)  	j=right;  	i=left;  	temp=a[left];  	                                 	if(left>right) return;  	int i,j,t,temp;  {  void QuickSortSecond(int left,int right,int a[NODENUM])   } 	return i; 	a[i]=temp;      a[left]=a[i];  	} 		} 			a[j]=t;  			a[i]=a[j];  			t=a[i];  		{  		if(i<j)  		while(a[i]<=temp && i<j) i++;  		while(a[j]>=temp && i<j) j--;  	{  	while(i!=j)  	j=right;  	i=left;  	temp=a[left];  	                                 	if(left>right) return;  	int i,j,t,temp;  {  int QuickSortFirst(int left,int right,int a[NODENUM])   }     fclose(fp);     printf("\n");     }                              }                 p=strtok(NULL," ");                 i++;                 c[i] = atoi(p);             {             while (p)             p=strtok(str," ");         if (fgets(str,sizeof(str),fp)==NULL) break ;         char *p;         char str[1024];     {     while(!feof(fp))         }         printf("open file error\n");     {     if (fp == NULL)     fp=fopen(contents,"r");     //begin to read file       FILE *fp;     int j;     int i = 0; void ReadFile(char *contents, int c[NODENUM]){  volatile int FinalArray[NODENUM+128]; volatile int InputArray[NODENUM];  extern void MTA_printresult();   #define LOCALNUM 250 #define NODENUM 500 #define INF 20000  #define cmp1_7 0x1ff008000 #define cmp1_6 0x1ff007000 #define cmp1_5 0x1ff006000 #define cmp1_4 0x1ff005000 #define cmp1_3 0x1ff004000 #define cmp1_2 0x1ff003000 #define cmp1_1 0x1ff002000 #define cmp1_0 0x1ff001000  #define cmp0_6 0x11fde6f50 #define cmp0_5 0x1ff000800 #define cmp0_4 0x1ff000400 #define cmp0_3 0x1ff000300 #define cmp0_2 0x1ff000200 #define cmp0_1 0x1ff000100 #define cmp0_0 0x1ff000000  volatile int CountLock = 0; #define NPROC 16  #include "stdint.h" #include "barrier.h" #include "stdio.h" #define global ad  
  �
     0       ]  .      �  �  �  �  �  �  I  )    �  �  �  �  �  |  {  j  7    �  �  �  �  �  �  w  s  p  o  Y  &  �  �  �  �  �  |  W  D  /    �
  �
  �
  �
  z
  y
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        } 	while(1); 	MTA_Stats(0);     //        MTA_tot} 	while(1); 	MTA_Stats(0);     //       } 	while(1); 	MTA_Stats(0); } 	while(1); 	MTA_Stats(0);     //        MTA_total_sim_cycle;     //if(my_id == 0) 	MTA_Bar_Stats(0); 	barrier(MTA_getthreadID() , NPROC); 	MTA_Bar_Stats(1);      }*/             fflush(stdout);             printf("The final sim-cycle is:%llu\n",finalSimCycle);             finalSimCycle = MTA_printresult();             printf("Print the final sim_cycle\n");     /*if(my_id == 0){  	} 		} 			WriteFile("./output.txt",FinalArray,NODENUM);             fflush(stdout); 			printf("The results is:\n"); 	if(my_id == 1){      }             MTA_printresult();             fflush(stdout);             printf("Print the final sim_cycle\n"); 	if(my_id == 0){  		MTA_Bar_Stats(0); 		barrier(MTA_getthreadID() , NPROC); 		MTA_Bar_Stats(1);          } 			MergeSort(FinalArray,0,LOCALNUM-1,NODENUM);             ReceiveData(FinalArray);             fflush(stdout);                 printf("I receive the data beginning...\n");              WaitTime(999);            if(my_id == 0){  		MTA_Bar_Stats(0); 		barrier(MTA_getthreadID() , NPROC); 		MTA_Bar_Stats(1);         }             fflush(stdout);             printf("This is the 64th loop\n"); 			MergeSort(FinalArray,my_id*(64*eachCoreNum),my_id*(64*eachCoreNum)+((((my_id+1)*64*eachCoreNum) -1)-my_id*(64*eachCoreNum))/2,((my_id+1)*(64*eachCoreNum)) -1); 